module MemoriaInstrucoes(Endereco,Clock,Instrucao);
	input [31:0] Endereco;
	input Clock;
	output [31:0] Instrucao;
	
	reg[31:0] Memory[255:0];
	integer F = 0;
	
	
	always @(posedge Clock)
	begin
	
		// Codigo	
		if(F == 0)
		begin
Memory[ 0] = 32'B00001000000000010000000000011010; // addi	$ra $zero 26
Memory[ 1] = 32'B00001000000111110000000001001100; // addi	$sp $zero 76
Memory[ 2] = 32'B00010100000000000000000001100101; // jump	main
Memory[ 3] = 32'B00110000000000000000000000000000; // nop	minloc
Memory[ 4] = 32'B00011100000000100000000000001010; // sw	$a0 10($zero)
Memory[ 5] = 32'B00011100000000110000000000001011; // sw	$a1 11($zero)
Memory[ 6] = 32'B00011100000001000000000000001100; // sw	$a2 12($zero)
Memory[ 7] = 32'B00011000000101010000000000001011; // lw	$s1 11($zero)
Memory[ 8] = 32'B00011100000101010000000000001111; // sw	$s1 15($zero)
Memory[ 9] = 32'B00011000000101010000000000001011; // lw	$s1 11($zero)
Memory[10] = 32'B00011000000101000000000000001010; // lw	$s0 10($zero)
Memory[11] = 32'B00000010100101011010000000000000; // add	$s0 $s0 $s1
Memory[12] = 32'B00011010100010000000000000000000; // lw	$t0 0($s0)
Memory[13] = 32'B00011100000010000000000000001110; // sw	$t0 14($zero)
Memory[14] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
Memory[15] = 32'B00011000000101000000000000001011; // lw	$s0 11($zero)
Memory[16] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
Memory[17] = 32'B00011100000010010000000000001101; // sw	$t1 13($zero)
Memory[18] = 32'B00110000000000000000000000000000; // nop	L0
Memory[19] = 32'B00011000000101000000000000001101; // lw	$s0 13($zero)
Memory[20] = 32'B00011000000101010000000000001100; // lw	$s1 12($zero)
Memory[21] = 32'B00010010100101010100000000000000; // slt	$t0 $s0 $s1
Memory[22] = 32'B00101001000000000000000000101101; // beq	$t0 0 L1
Memory[23] = 32'B00011000000101010000000000001101; // lw	$s1 13($zero)
Memory[24] = 32'B00011000000101000000000000001010; // lw	$s0 10($zero)
Memory[25] = 32'B00000010100101011010000000000000; // add	$s0 $s0 $s1
Memory[26] = 32'B00011010100010010000000000000000; // lw	$t1 0($s0)
Memory[27] = 32'B00011000000101010000000000001110; // lw	$s1 14($zero)
Memory[28] = 32'B00010001001101010101000000000000; // slt	$t2 $t1 $s1
Memory[29] = 32'B00101001010000000000000000100110; // beq	$t2 0 L2
Memory[30] = 32'B00011000000101010000000000001101; // lw	$s1 13($zero)
Memory[31] = 32'B00011000000101000000000000001010; // lw	$s0 10($zero)
Memory[32] = 32'B00000010100101011010000000000000; // add	$s0 $s0 $s1
Memory[33] = 32'B00011010100010110000000000000000; // lw	$t3 0($s0)
Memory[34] = 32'B00011100000010110000000000001110; // sw	$t3 14($zero)
Memory[35] = 32'B00011000000101010000000000001101; // lw	$s1 13($zero)
Memory[36] = 32'B00011100000101010000000000001111; // sw	$s1 15($zero)
Memory[37] = 32'B00010100000000000000000000100111; // jump	L3
Memory[38] = 32'B00110000000000000000000000000000; // nop	L2
Memory[39] = 32'B00110000000000000000000000000000; // nop	L3
Memory[40] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
Memory[41] = 32'B00011000000101000000000000001101; // lw	$s0 13($zero)
Memory[42] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
Memory[43] = 32'B00011100000010010000000000001101; // sw	$t1 13($zero)
Memory[44] = 32'B00010100000000000000000000010010; // jump	L0
Memory[45] = 32'B00110000000000000000000000000000; // nop	L1
Memory[46] = 32'B00011000000101010000000000001111; // lw	$s1 15($zero)
Memory[47] = 32'B00001110101111100000000000000000; // move	$v0 $s1 
Memory[48] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
Memory[49] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
Memory[50] = 32'B01001110100000000000000000000000; // jr	$s0  
Memory[51] = 32'B00110000000000000000000000000000; // nop	sort
Memory[52] = 32'B00011100000000100000000000010000; // sw	$a0 16($zero)
Memory[53] = 32'B00011100000000110000000000010001; // sw	$a1 17($zero)
Memory[54] = 32'B00011100000001000000000000010010; // sw	$a2 18($zero)
Memory[55] = 32'B00011000000101010000000000010001; // lw	$s1 17($zero)
Memory[56] = 32'B00011100000101010000000000010011; // sw	$s1 19($zero)
Memory[57] = 32'B00110000000000000000000000000000; // nop	L4
Memory[58] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
Memory[59] = 32'B00011000000101000000000000010010; // lw	$s0 18($zero)
Memory[60] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
Memory[61] = 32'B00011000000101000000000000010011; // lw	$s0 19($zero)
Memory[62] = 32'B00010010100010010101000000000000; // slt	$t2 $s0 $t1
Memory[63] = 32'B00101001010000000000000001100001; // beq	$t2 0 L5
Memory[64] = 32'B00011000000000100000000000010000; // lw	$a0 16($zero)
Memory[65] = 32'B00011000000101010000000000010011; // lw	$s1 19($zero)
Memory[66] = 32'B00001110101000110000000000000000; // move	$a1 $s1 
Memory[67] = 32'B00011000000101010000000000010010; // lw	$s1 18($zero)
Memory[68] = 32'B00001110101001000000000000000000; // move	$a2 $s1 
Memory[69] = 32'B00001000000101000000000001001001; // addi	$s0 $zero 73
Memory[70] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
Memory[71] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
Memory[72] = 32'B00010100000000000000000000000011; // jump	minloc
Memory[73] = 32'B00011100000111100000000000010100; // sw	$v0 20($zero)
Memory[74] = 32'B00011000000101010000000000010100; // lw	$s1 20($zero)
Memory[75] = 32'B00011000000101000000000000010000; // lw	$s0 16($zero)
Memory[76] = 32'B00000010100101011010000000000000; // add	$s0 $s0 $s1
Memory[77] = 32'B00011010100010000000000000000000; // lw	$t0 0($s0)
Memory[78] = 32'B00011100000010000000000000010101; // sw	$t0 21($zero)
Memory[79] = 32'B00011000000101010000000000010011; // lw	$s1 19($zero)
Memory[80] = 32'B00011000000101000000000000010000; // lw	$s0 16($zero)
Memory[81] = 32'B00000010100101011010000000000000; // add	$s0 $s0 $s1
Memory[82] = 32'B00011010100010000000000000000000; // lw	$t0 0($s0)
Memory[83] = 32'B00011000000101000000000000010000; // lw	$s0 16($zero)
Memory[84] = 32'B00011000000101010000000000010100; // lw	$s1 20($zero)
Memory[85] = 32'B00000010101101000100100000000000; // add	$t1 $s0 $s1
Memory[86] = 32'B00011101001010000000000000000000; // sw	$t0 0($t1)
Memory[87] = 32'B00011000000101000000000000010000; // lw	$s0 16($zero)
Memory[88] = 32'B00011000000101010000000000010011; // lw	$s1 19($zero)
Memory[89] = 32'B00000010101101000100000000000000; // add	$t0 $s0 $s1
Memory[90] = 32'B00011000000101010000000000010101; // lw	$s1 21($zero)
Memory[91] = 32'B00011101000101010000000000000000; // sw	$s1 0($t0)
Memory[92] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
Memory[93] = 32'B00011000000101000000000000010011; // lw	$s0 19($zero)
Memory[94] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
Memory[95] = 32'B00011100000010010000000000010011; // sw	$t1 19($zero)
Memory[96] = 32'B00010100000000000000000000111001; // jump	L4
Memory[97] = 32'B00110000000000000000000000000000; // nop	L5
Memory[98] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
Memory[99] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
Memory[100] = 32'B01001110100000000000000000000000; // jr	$s0  
Memory[101] = 32'B00110000000000000000000000000000; // nop	main
Memory[102] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
Memory[103] = 32'B00011100000010000000000000010111; // sw	$t0 23($zero)
Memory[104] = 32'B00110000000000000000000000000000; // nop	L6
Memory[105] = 32'B00001000000010000000000000001010; // addi	$t0 $zero 10
Memory[106] = 32'B00011000000101000000000000010111; // lw	$s0 23($zero)
Memory[107] = 32'B00010010100010000100100000000000; // slt	$t1 $s0 $t0
Memory[108] = 32'B00101001001000000000000001111010; // beq	$t1 0 L7
Memory[109] = 32'B00001000000010100000000000010100; // addi	$t2 $zero 20
Memory[110] = 32'B00001000000010110000000000000010; // addi	$t3 $zero 2
Memory[111] = 32'B00011000000101010000000000010111; // lw	$s1 23($zero)
Memory[112] = 32'B00000001011101010110000000000010; // mult	$t4 $t3 $s1
Memory[113] = 32'B00000001010011000110100000000001; // sub	$t5 $t2 $t4
Memory[114] = 32'B00011000000101010000000000010111; // lw	$s1 23($zero)
Memory[115] = 32'B00001010101011100000000000000000; // addi	$t6 $s1 0
Memory[116] = 32'B00011101110011010000000000000000; // sw	$t5 0($t6)
Memory[117] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
Memory[118] = 32'B00011000000101000000000000010111; // lw	$s0 23($zero)
Memory[119] = 32'B00000001000101000100100000000000; // add	$t1 $s0 $t0
Memory[120] = 32'B00011100000010010000000000010111; // sw	$t1 23($zero)
Memory[121] = 32'B00010100000000000000000001101000; // jump	L6
Memory[122] = 32'B00110000000000000000000000000000; // nop	L7
Memory[123] = 32'B00001000000000100000000000000000; // addi	$a0 $zero 0
Memory[124] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
Memory[125] = 32'B00001101000000110000000000000000; // move	$a1 $t0 
Memory[126] = 32'B00001000000010010000000000001010; // addi	$t1 $zero 10
Memory[127] = 32'B00001101001001000000000000000000; // move	$a2 $t1 
Memory[128] = 32'B00001000000101000000000010000100; // addi	$s0 $zero 132
Memory[129] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
Memory[130] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
Memory[131] = 32'B00010100000000000000000000110011; // jump	sort
Memory[132] = 32'B00001000000010100000000000000000; // addi	$t2 $zero 0
Memory[133] = 32'B00011100000010100000000000010111; // sw	$t2 23($zero)
Memory[134] = 32'B00110000000000000000000000000000; // nop	L8
Memory[135] = 32'B00001000000010000000000000001010; // addi	$t0 $zero 10
Memory[136] = 32'B00011000000101000000000000010111; // lw	$s0 23($zero)
Memory[137] = 32'B00010010100010000100100000000000; // slt	$t1 $s0 $t0
Memory[138] = 32'B00101001001000000000000010010100; // beq	$t1 0 L9
Memory[139] = 32'B00011000000101010000000000010111; // lw	$s1 23($zero)
Memory[140] = 32'B00011010101010100000000000000000; // lw	$t2 0($s1)
Memory[141] = 32'B00001101010000100000000000000000; // move	$a0 $t2 
Memory[142] = 32'B00100100010000000000000000000000; // out	$a0  
Memory[143] = 32'B00001000000010110000000000000001; // addi	$t3 $zero 1
Memory[144] = 32'B00011000000101000000000000010111; // lw	$s0 23($zero)
Memory[145] = 32'B00000001011101000110000000000000; // add	$t4 $s0 $t3
Memory[146] = 32'B00011100000011000000000000010111; // sw	$t4 23($zero)
Memory[147] = 32'B00010100000000000000000010000110; // jump	L8
Memory[148] = 32'B00110000000000000000000000000000; // nop	L9
Memory[149] = 32'B00010100000000000000000010010101; // halt	    
		F = 1;
		end
		///////////////////////////////////
	end
	
	assign Instrucao = Memory[Endereco];
	
endmodule
