module MemoriaInstrucoes(Endereco,Clock,Instrucao);
	input [31:0] Endereco;
	input Clock;
	output [31:0] Instrucao;
	
	reg[31:0] Memory[122:0];
	integer F = 0;
	
	
	always @(posedge Clock)
	begin
	
		// Codigo	
		if(F == 0)
		begin
		Memory[ 0] = 32'B00001000000000010000000000001001; // addi	$ra $zero 9
		Memory[ 1] = 32'B00001000000111110000000000111011; // addi	$sp $zero 59
		Memory[ 2] = 32'B00010100000000000000000000101000; // jump	main
		Memory[ 3] = 32'B00110000000000000000000000000000; // nop	Combinatoria
		Memory[ 4] = 32'B00011100000000100000000000000000; // sw	$a0 0($zero)
		Memory[ 5] = 32'B00011100000000110000000000000001; // sw	$a1 1($zero)
		Memory[ 6] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		Memory[ 7] = 32'B00011100000010000000000000000010; // sw	$t0 2($zero)
		Memory[ 8] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		Memory[ 9] = 32'B00011100000010000000000000000011; // sw	$t0 3($zero)
		Memory[10] = 32'B00110000000000000000000000000000; // nop	L0
		Memory[11] = 32'B00001000000010000000000000000000; // addi	$t0 $zero 0
		Memory[12] = 32'B00011000000101000000000000000001; // lw	$s0 1($zero)
		Memory[13] = 32'B00111110100010000100100000000000; // sbt	$t1 $s0 $t0
		Memory[14] = 32'B00101001001000000000000000100000; // beq	$t1 0 L1
		Memory[15] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		Memory[16] = 32'B00011000000101010000000000000000; // lw	$s1 0($zero)
		Memory[17] = 32'B00000010100101010101000000000010; // mult	$t2 $s0 $s1
		Memory[18] = 32'B00011100000010100000000000000010; // sw	$t2 2($zero)
		Memory[19] = 32'B00011000000101000000000000000011; // lw	$s0 3($zero)
		Memory[20] = 32'B00011000000101010000000000000001; // lw	$s1 1($zero)
		Memory[21] = 32'B00000010100101010100000000000010; // mult	$t0 $s0 $s1
		Memory[22] = 32'B00011100000010000000000000000011; // sw	$t0 3($zero)
		Memory[23] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		Memory[24] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
		Memory[25] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
		Memory[26] = 32'B00011100000010010000000000000000; // sw	$t1 0($zero)
		Memory[27] = 32'B00001000000010000000000000000001; // addi	$t0 $zero 1
		Memory[28] = 32'B00011000000101000000000000000001; // lw	$s0 1($zero)
		Memory[29] = 32'B00000010100010000100100000000001; // sub	$t1 $s0 $t0
		Memory[30] = 32'B00011100000010010000000000000001; // sw	$t1 1($zero)
		Memory[31] = 32'B00010100000000000000000000001010; // jump	L0
		Memory[32] = 32'B00110000000000000000000000000000; // nop	L1
		Memory[33] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
		Memory[34] = 32'B00011000000101010000000000000011; // lw	$s1 3($zero)
		Memory[35] = 32'B00000010100101010100000000000011; // div	$t0 $s0 $s1
		Memory[36] = 32'B00001101000111100000000000000000; // move	$v0 $t0 
		Memory[37] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
		Memory[38] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
		Memory[39] = 32'B01001110100000000000000000000000; // jr	$s0  
		Memory[40] = 32'B00110000000000000000000000000000; // nop	main
		Memory[41] = 32'B00100000010000100000000000000000; // in	$a0  
		Memory[42] = 32'B00011100000000100000000000000100; // sw	$a0 4($zero)
		Memory[43] = 32'B00100000010000100000000000000000; // in	$a0  
		Memory[44] = 32'B00011100000000100000000000000101; // sw	$a0 5($zero)
		Memory[45] = 32'B00011000000101010000000000000100; // lw	$s1 4($zero)
		Memory[46] = 32'B00001110101000100000000000000000; // move	$a0 $s1 
		Memory[47] = 32'B00011000000101010000000000000101; // lw	$s1 5($zero)
		Memory[48] = 32'B00001110101000110000000000000000; // move	$a1 $s1 
		Memory[49] = 32'B00001000000101000000000000110101; // addi	$s0 $zero 53
		Memory[50] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
		Memory[51] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
		Memory[52] = 32'B00010100000000000000000000000011; // jump	Combinatoria
		Memory[53] = 32'B00001111110001000000000000000000; // move	$a2 $v0 
		Memory[54] = 32'B00100100100000000000000000000000; // out	$a2  
		Memory[55] = 32'B00010100000000000000000000110111; // halt	   	         	                        
		F = 1;
		end
		///////////////////////////////////
	end
	
	assign Instrucao = Memory[Endereco];
	
endmodule
