module MemoriaInstrucoes(Endereco,Clock,Instrucao);
	input [31:0] Endereco;
	input Clock;
	output [31:0] Instrucao;
	
	reg[31:0] Memory[52:0];
	integer F = 0;
	
	
	always @(posedge Clock)
	begin
	
		// Codigo	
		if(F == 0)
		begin	
		
Memory[ 0] = 32'B00001000000000010000000000110010; // addi	$ra $zero 50
Memory[ 1] = 32'B00001000000111110000000001001011; // addi	$sp $zero 75
Memory[ 2] = 32'B00010100000000000000000000011001; // jump	main
Memory[ 3] = 32'B00110000000000000000000000000000; // nop	PreencherVetor
Memory[ 4] = 32'B00011100000000100000000000000000; // sw	$a0 0($zero)
Memory[ 5] = 32'B00011100000000110000000000000001; // sw	$a1 1($zero)
Memory[ 6] = 32'B00001000000001110000000000000000; // addi	$t0 $zero 0
Memory[ 7] = 32'B00011100000001110000000000000010; // sw	$t0 2($zero)
Memory[ 8] = 32'B00110000000000000000000000000000; // nop	L0
Memory[ 9] = 32'B00011000000101000000000000000010; // lw	$s0 2($zero)
Memory[10] = 32'B00011000000101010000000000000001; // lw	$s1 1($zero)
Memory[11] = 32'B00010010100101010011100000000000; // slt	$t0 $s0 $s1
Memory[12] = 32'B00101000111000000000000000010101; // beq	$t0 0 L1
Memory[13] = 32'B00001000000010000000000000000010; // addi	$t1 $zero 2
Memory[14] = 32'B00011000000101010000000000000010; // lw	$s1 2($zero)
Memory[15] = 32'B00000001000101010100100000000010; // mult	$t2 $t1 $s1
Memory[16] = 32'B00011000000101000000000000000000; // lw	$s0 0($zero)
Memory[17] = 32'B00011000000101010000000000000010; // lw	$s1 2($zero)
Memory[18] = 32'B00000010101101000101000000000000; // add	$t3 $s0 $s1
Memory[19] = 32'B00011101010010010000000000000000; // sw	$t2 0($t3)
Memory[20] = 32'B00010100000000000000000000001000; // jump	L0
Memory[21] = 32'B00110000000000000000000000000000; // nop	L1
Memory[22] = 32'B01010000001000010000000000000001; // subi	$ra $ra 1
Memory[23] = 32'B00011000001101000000000000000000; // lw	$s0 0($ra)
Memory[24] = 32'B01001110100000000000000000000000; // jr	$s0  
Memory[25] = 32'B00110000000000000000000000000000; // nop	main
Memory[26] = 32'B00001000000001110000000000001111; // addi	$t0 $zero 15
Memory[27] = 32'B00011100000001110000000000000100; // sw	$t0 4($zero)
Memory[28] = 32'B00001000000000100000000000000101; // addi	$a0 $zero 5
Memory[29] = 32'B00011000000101010000000000000100; // lw	$s1 4($zero)
Memory[30] = 32'B00001110101000110000000000000000; // move	$a1 $s1 
Memory[31] = 32'B00001000000101000000000000100011; // addi	$s0 $zero 35
Memory[32] = 32'B00011100001101000000000000000000; // sw	$s0 0($ra)
Memory[33] = 32'B00001000001000010000000000000001; // addi	$ra $ra 1
Memory[34] = 32'B00010100000000000000000000000011; // jump	PreencherVetor
Memory[35] = 32'B00001000000001110000000000000000; // addi	$t0 $zero 0
Memory[36] = 32'B00011100000001110000000000000011; // sw	$t0 3($zero)
Memory[37] = 32'B00110000000000000000000000000000; // nop	L2
Memory[38] = 32'B00011000000101000000000000000011; // lw	$s0 3($zero)
Memory[39] = 32'B00011000000101010000000000000100; // lw	$s1 4($zero)
Memory[40] = 32'B00010010100101010011100000000000; // slt	$t0 $s0 $s1
Memory[41] = 32'B00101000111000000000000000110011; // beq	$t0 0 L3
Memory[42] = 32'B00011000000101010000000000000011; // lw	$s1 3($zero)
Memory[43] = 32'B00011010101010000000000000000101; // lw	$t1 5($s1)
Memory[44] = 32'B00001101000000100000000000000000; // move	$a0 $t1 
Memory[45] = 32'B00100100010000000000000000000000; // out	$a0  
Memory[46] = 32'B00001000000010010000000000000001; // addi	$t2 $zero 1
Memory[47] = 32'B00011000000101000000000000000011; // lw	$s0 3($zero)
Memory[48] = 32'B00000001001101000101000000000000; // add	$t3 $s0 $t2
Memory[49] = 32'B00011100000010100000000000000011; // sw	$t3 3($zero)
Memory[50] = 32'B00010100000000000000000000100101; // jump	L2
Memory[51] = 32'B00110000000000000000000000000000; // nop	L3
Memory[52] = 32'B00010100000000000000000000110100; // halt	  

		F = 1;
		end
		///////////////////////////////////
	end
	
	assign Instrucao = Memory[Endereco];
	
endmodule
